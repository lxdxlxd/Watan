6
0 0 0 1 0 g 0 0 c 0 1 50 1 
0 0 0 1 0 g 0 0 c 4 1 46 1 
0 0 1 0 0 g 0 0 c 10 1 41 1 
0 0 1 0 0 g 0 0 c 17 1 29 1 
1 10 3 8 3 6 0 8 2 3 2 4 4 10 0 9 2 11 1 6 1 2 0 5 5 7 0 5 4 11 1 3 2 12 3 4 4 9 
14